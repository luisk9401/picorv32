// Environment for simpleuart
class simpleuart_env extends uvm_env;
    simpleuart_agent agent;
    `uvm_component_utils(simpleuart_env)
endclass
