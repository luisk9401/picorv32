package picorv32_axi_adapter_types;

    typedef enum {READ, WRITE, RESET} a_tran_type; 

endpackage : picorv32_axi_adapter_types
