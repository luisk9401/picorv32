package sequences_pkg;

   import uvm_pkg::*;
   import picorv32_axi_adapter_pkg::*;
   `include "uvm_macros.svh"
   `include "sequences/basic_read_write_sequence.sv"
   //`include "sequences/invalid_state_sequence.sv"
   //`include "sequences/simultaneous_read_write_sequence.sv"
endpackage : sequences_pkg
