// Interface for simpleuart
interface simpleuart_if(input logic clk, input logic resetn);
    logic [7:0] data;
endinterface
