// Environment for spimemio
class spimemio_env extends uvm_env;
    spimemio_agent agent;
    `uvm_component_utils(spimemio_env)
endclass
