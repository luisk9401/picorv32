package pcpi_div_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "pcpi_div_txn.sv"
    `include "pcpi_div_sqr.sv"
    `include "pcpi_div_mon.sv"
    `include "pcpi_div_drv.sv"
    //`include "pcpi_div_adapter.sv"
    `include "pcpi_div_agent.sv"
endpackage
