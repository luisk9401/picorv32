//===============================================================
// Top HVL for Full Chip Environment
//===============================================================
module top_hvl;
    import uvm_pkg::*;
    import fullchip_pkg::*;
    initial begin
        run_test();
    end
endmodule
